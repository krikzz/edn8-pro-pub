

	`define SST_ON	//save state
	`define CCO_ON	//cheats codes engine
	`define SND_ON	//expansion sound if any exists
